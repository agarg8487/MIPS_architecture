/* 
Authors : Aditya Terkar, 16EC01003, IIT Bhubaneswar
Aim : 
*/
//////////////////////////////////////////////////////////////////////////////////////////
//project includes
/////////////////////////////////////////////////////////////////////////////////////////

module mod_write_data_mux ( 
                            //input ports
                            input [31 : 0] ext_mem_data,
                            input [31 : 0] alu_data,
                            input mem_to_reg,
                            
                            //output ports
                            output wire [31 : 0] write_data
                          );
//----------------------------parameters---------------------------------
//-----------------------------------------------------------------------
//-------------------------module instantiation--------------------------
//-----------------------------------------------------------------------
//-------------------------hardware action-------------------------------
    assign write_data = (mem_to_reg) ? ext_mem_data : alu_data;
//-----------------------------------------------------------------------
//----------------------functions and tasks------------------------------
//-----------------------------------------------------------------------
endmodule