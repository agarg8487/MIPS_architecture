/* 
Authors : Adtiya Terkar, 16EC01003, IIT Bhubaneswar
Aim : A instruction provider
*/ 
//////////////////////////////////////////////////////////////////////////////////////////
//project includes
/////////////////////////////////////////////////////////////////////////////////////////
module mod_instruction_mem_rom (
    //input ports
    input [29 : 0] address,
    //output ports
    output reg [31 : 0] instruction,
    output wire mem_end);

//-------------------------hardware action-------------------------------
    always @(*) begin
        case (address)
            0 : instruction = 32'b00000100000000000000000000000001;
            1 : instruction = 32'b00000100000000010000000000000010;
            2 : instruction = 32'b00000100000000100000000000000011;
            3 : instruction = 32'b00000100000000110000000000000100;
            4 : instruction = 32'b00000100000001000000000000000100;
            5 : instruction = 32'b00010000011001001111111111111110;
            6 : instruction = 32'b00000100000001010000000000000110;
            7 : instruction = 32'b00000100000001100000000000000111;
            8 : instruction = 32'b00000100000001110000000000001000;
            9 : instruction = 32'b00000100000010000000000000001001;
            10 : instruction = 32'b00000100000010010000000000001010;
            11 : instruction = 32'b00000100000010100000000000001011;
            12 : instruction = 32'b00000100000010110000000000001100;
            13 : instruction = 32'b00000100000011000000000000001101;
            14 : instruction = 32'b00000100000011010000000000001110;
            15 : instruction = 32'b00000100000011100000000000001111;
            16 : instruction = 32'b00000100000011110000000000010000;
            17 : instruction = 32'b00000100000100000000000000010001;
            18 : instruction = 32'b00000100000100010000000000010010;
            19 : instruction = 32'b00000100000100100000000000010011;
            20 : instruction = 32'b00000100000100110000000000010100;
            21 : instruction = 32'b00000100000101000000000000010101;
            22 : instruction = 32'b00000100000101010000000000010110;
            23 : instruction = 32'b00000100000101100000000000010111;
            24 : instruction = 32'b00000100000101110000000000011000;
            25 : instruction = 32'b00000100000110000000000000011001;
            26 : instruction = 32'b00000100000110010000000000011010;
            27 : instruction = 32'b00000100000110100000000000011011;
            28 : instruction = 32'b00000100000110110000000000011100;
            29 : instruction = 32'b00000100000111000000000000011101;
            30 : instruction = 32'b00000100000111010000000000011110;
            31 : instruction = 32'b00000100000111100000000000011111;
            32 : instruction = 32'b00000100000111110000000000100000;
            33 : instruction = 32'b00000000010000000000100000100000;
            34 : instruction = 32'b00000000000000000001100000100000;
            default : instruction = 0;
        endcase
    end
    assign mem_end = (address > 34) ? 1'b1 : 1'b0;//-----------------------------------------------------------------------
endmodule
