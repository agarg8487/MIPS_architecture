/* 
Authors : Adtiya Terkar, 16EC01003, IIT Bhubaneswar
Aim : 
*/
//////////////////////////////////////////////////////////////////////////////////////////
//project includes
/////////////////////////////////////////////////////////////////////////////////////////

module mod_pc_mux (input mux_control,
                            input [31 : 0] pc_plus_4,
                            input [31 : 0] branch_address,
                            output [31 : 0] next_address
                           );
//----------------------------parameters----------------------------------

//-----------------------------------------------------------------------
//-------------------------module instantiation--------------------------
//-----------------------------------------------------------------------
//-------------------------hardware action-------------------------------
//-----------------------------------------------------------------------
//----------------------functions and tasks------------------------------
//-----------------------------------------------------------------------
endmodule