/* 
Authors : Adtiya Terkar, 16EC01003, IIT Bhubaneswar
Aim : A instruction provider
*/ 
//////////////////////////////////////////////////////////////////////////////////////////
//project includes
/////////////////////////////////////////////////////////////////////////////////////////
module mod_instruction_mem_rom (
    //input ports
    input [29 : 0] address,
    //output ports
    output reg [31 : 0] instruction,
    output wire mem_end);

//-------------------------hardware action-------------------------------
    always @(*) begin
        case (address)
            0 : instruction = 32'b00100000000000010000000000000001;
            1 : instruction = 32'b00000000000000010001000000100000;
            2 : instruction = 32'b00001100000000010000000000000001;
            3 : instruction = 32'b00001100000000010000000000000010;
            4 : instruction = 32'b00100000000001010000000000010010;
            5 : instruction = 32'b00100000000001100000000000000001;
            6 : instruction = 32'b00100000000001110000000000000010;
            7 : instruction = 32'b00000000010000010001100000100000;
            8 : instruction = 32'b00100000111001110000000000000001;
            9 : instruction = 32'b00001100111000110000000000000000;
            10 : instruction = 32'b00000000000000100000100000100000;
            11 : instruction = 32'b00000000000000110001000000100000;
            12 : instruction = 32'b00000000101001100010100000100010;
            13 : instruction = 32'b00010000101000000000000000000001;
            14 : instruction = 32'b00001000000000000000000000000111;
            15 : instruction = 32'b00100000000010000011001101110010;
            16 : instruction = 32'b00100000111001110000000000000001;
            17 : instruction = 32'b00001100111010000000000000000000;
            18 : instruction = 32'b00100000000010010000000000000000;
            19 : instruction = 32'b00100000000010100000000000000000;
            20 : instruction = 32'b00000001000010100100100000101010;
            21 : instruction = 32'b00100000111001110000000000000001;
            22 : instruction = 32'b00001100111010010000000000000000;
            default : instruction = 0;
        endcase
    end
    assign mem_end = (address > 22) ? 1'b1 : 1'b0;//-----------------------------------------------------------------------
endmodule
